// IntegracaoPlatformDesigner.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module IntegracaoPlatformDesigner (
		input  wire        clk_clk,                       //                     clk.clk
		input  wire        reset_reset_n,                 //                   reset.reset_n
		input  wire        sram_conduit_cdt_write,        //            sram_conduit.cdt_write
		input  wire        sram_conduit_cdt_chipselect,   //                        .cdt_chipselect
		input  wire        sram_conduit_cdt_outputenable, //                        .cdt_outputenable
		input  wire [19:0] sram_conduit_cdt_address,      //                        .cdt_address
		inout  wire [15:0] sram_conduit_cdt_data_io,      //                        .cdt_data_io
		input  wire [1:0]  sram_conduit_cdt_byteenable,   //                        .cdt_byteenable
		inout  wire [15:0] sram_controller_conduit_DQ,    // sram_controller_conduit.DQ
		output wire [19:0] sram_controller_conduit_ADDR,  //                        .ADDR
		output wire        sram_controller_conduit_LB_N,  //                        .LB_N
		output wire        sram_controller_conduit_UB_N,  //                        .UB_N
		output wire        sram_controller_conduit_CE_N,  //                        .CE_N
		output wire        sram_controller_conduit_OE_N,  //                        .OE_N
		output wire        sram_controller_conduit_WE_N,  //                        .WE_N
		output wire        vga_conduit_CLK,               //             vga_conduit.CLK
		output wire        vga_conduit_HS,                //                        .HS
		output wire        vga_conduit_VS,                //                        .VS
		output wire        vga_conduit_BLANK,             //                        .BLANK
		output wire        vga_conduit_SYNC,              //                        .SYNC
		output wire [7:0]  vga_conduit_R,                 //                        .R
		output wire [7:0]  vga_conduit_G,                 //                        .G
		output wire [7:0]  vga_conduit_B                  //                        .B
	);

	wire         grayscale_converter_avalon_csc_source_valid;                       // grayscale_converter:stream_out_valid -> edge_detector:in_valid
	wire   [7:0] grayscale_converter_avalon_csc_source_data;                        // grayscale_converter:stream_out_data -> edge_detector:in_data
	wire         grayscale_converter_avalon_csc_source_ready;                       // edge_detector:in_ready -> grayscale_converter:stream_out_ready
	wire         grayscale_converter_avalon_csc_source_startofpacket;               // grayscale_converter:stream_out_startofpacket -> edge_detector:in_startofpacket
	wire         grayscale_converter_avalon_csc_source_endofpacket;                 // grayscale_converter:stream_out_endofpacket -> edge_detector:in_endofpacket
	wire         dual_clock_buffer_avalon_dc_buffer_source_valid;                   // dual_clock_buffer:stream_out_valid -> vga_controller:valid
	wire  [29:0] dual_clock_buffer_avalon_dc_buffer_source_data;                    // dual_clock_buffer:stream_out_data -> vga_controller:data
	wire         dual_clock_buffer_avalon_dc_buffer_source_ready;                   // vga_controller:ready -> dual_clock_buffer:stream_out_ready
	wire         dual_clock_buffer_avalon_dc_buffer_source_startofpacket;           // dual_clock_buffer:stream_out_startofpacket -> vga_controller:startofpacket
	wire         dual_clock_buffer_avalon_dc_buffer_source_endofpacket;             // dual_clock_buffer:stream_out_endofpacket -> vga_controller:endofpacket
	wire         edge_detector_avalon_edge_detection_source_valid;                  // edge_detector:out_valid -> resample_1bit:stream_in_valid
	wire   [7:0] edge_detector_avalon_edge_detection_source_data;                   // edge_detector:out_data -> resample_1bit:stream_in_data
	wire         edge_detector_avalon_edge_detection_source_ready;                  // resample_1bit:stream_in_ready -> edge_detector:out_ready
	wire         edge_detector_avalon_edge_detection_source_startofpacket;          // edge_detector:out_startofpacket -> resample_1bit:stream_in_startofpacket
	wire         edge_detector_avalon_edge_detection_source_endofpacket;            // edge_detector:out_endofpacket -> resample_1bit:stream_in_endofpacket
	wire         pixel_buffer_avalon_pixel_source_valid;                            // pixel_buffer:stream_valid -> resample_24bit:stream_in_valid
	wire  [15:0] pixel_buffer_avalon_pixel_source_data;                             // pixel_buffer:stream_data -> resample_24bit:stream_in_data
	wire         pixel_buffer_avalon_pixel_source_ready;                            // resample_24bit:stream_in_ready -> pixel_buffer:stream_ready
	wire         pixel_buffer_avalon_pixel_source_startofpacket;                    // pixel_buffer:stream_startofpacket -> resample_24bit:stream_in_startofpacket
	wire         pixel_buffer_avalon_pixel_source_endofpacket;                      // pixel_buffer:stream_endofpacket -> resample_24bit:stream_in_endofpacket
	wire         resample_24bit_avalon_rgb_source_valid;                            // resample_24bit:stream_out_valid -> grayscale_converter:stream_in_valid
	wire  [23:0] resample_24bit_avalon_rgb_source_data;                             // resample_24bit:stream_out_data -> grayscale_converter:stream_in_data
	wire         resample_24bit_avalon_rgb_source_ready;                            // grayscale_converter:stream_in_ready -> resample_24bit:stream_out_ready
	wire         resample_24bit_avalon_rgb_source_startofpacket;                    // resample_24bit:stream_out_startofpacket -> grayscale_converter:stream_in_startofpacket
	wire         resample_24bit_avalon_rgb_source_endofpacket;                      // resample_24bit:stream_out_endofpacket -> grayscale_converter:stream_in_endofpacket
	wire         resample_1bit_avalon_rgb_source_valid;                             // resample_1bit:stream_out_valid -> vga_resample:stream_in_valid
	wire         resample_1bit_avalon_rgb_source_data;                              // resample_1bit:stream_out_data -> vga_resample:stream_in_data
	wire         resample_1bit_avalon_rgb_source_ready;                             // vga_resample:stream_in_ready -> resample_1bit:stream_out_ready
	wire         resample_1bit_avalon_rgb_source_startofpacket;                     // resample_1bit:stream_out_startofpacket -> vga_resample:stream_in_startofpacket
	wire         resample_1bit_avalon_rgb_source_endofpacket;                       // resample_1bit:stream_out_endofpacket -> vga_resample:stream_in_endofpacket
	wire         vga_resample_avalon_rgb_source_valid;                              // vga_resample:stream_out_valid -> scaler:stream_in_valid
	wire  [29:0] vga_resample_avalon_rgb_source_data;                               // vga_resample:stream_out_data -> scaler:stream_in_data
	wire         vga_resample_avalon_rgb_source_ready;                              // scaler:stream_in_ready -> vga_resample:stream_out_ready
	wire         vga_resample_avalon_rgb_source_startofpacket;                      // vga_resample:stream_out_startofpacket -> scaler:stream_in_startofpacket
	wire         vga_resample_avalon_rgb_source_endofpacket;                        // vga_resample:stream_out_endofpacket -> scaler:stream_in_endofpacket
	wire         scaler_avalon_scaler_source_valid;                                 // scaler:stream_out_valid -> dual_clock_buffer:stream_in_valid
	wire  [29:0] scaler_avalon_scaler_source_data;                                  // scaler:stream_out_data -> dual_clock_buffer:stream_in_data
	wire         scaler_avalon_scaler_source_ready;                                 // dual_clock_buffer:stream_in_ready -> scaler:stream_out_ready
	wire         scaler_avalon_scaler_source_startofpacket;                         // scaler:stream_out_startofpacket -> dual_clock_buffer:stream_in_startofpacket
	wire         scaler_avalon_scaler_source_endofpacket;                           // scaler:stream_out_endofpacket -> dual_clock_buffer:stream_in_endofpacket
	wire         pll_vga_vga_clk_clk;                                               // pll_vga:vga_clk_clk -> [dual_clock_buffer:clk_stream_out, rst_controller_001:clk, rst_controller_002:clk, vga_controller:clk]
	wire         pixel_buffer_avalon_pixel_dma_master_waitrequest;                  // mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_waitrequest -> pixel_buffer:master_waitrequest
	wire  [15:0] pixel_buffer_avalon_pixel_dma_master_readdata;                     // mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_readdata -> pixel_buffer:master_readdata
	wire  [31:0] pixel_buffer_avalon_pixel_dma_master_address;                      // pixel_buffer:master_address -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_address
	wire         pixel_buffer_avalon_pixel_dma_master_read;                         // pixel_buffer:master_read -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_read
	wire         pixel_buffer_avalon_pixel_dma_master_readdatavalid;                // mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_readdatavalid -> pixel_buffer:master_readdatavalid
	wire         pixel_buffer_avalon_pixel_dma_master_lock;                         // pixel_buffer:master_arbiterlock -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_lock
	wire  [31:0] nios_data_master_readdata;                                         // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                                      // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                                      // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [21:0] nios_data_master_address;                                          // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                                       // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                             // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                                            // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                        // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                                  // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                               // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [21:0] nios_instruction_master_address;                                   // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                                      // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire  [15:0] mm_interconnect_0_sram_controller_avalon_sram_slave_readdata;      // sram_controller:readdata -> mm_interconnect_0:sram_controller_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_controller_avalon_sram_slave_address;       // mm_interconnect_0:sram_controller_avalon_sram_slave_address -> sram_controller:address
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_read;          // mm_interconnect_0:sram_controller_avalon_sram_slave_read -> sram_controller:read
	wire   [1:0] mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable;    // mm_interconnect_0:sram_controller_avalon_sram_slave_byteenable -> sram_controller:byteenable
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid; // sram_controller:readdatavalid -> mm_interconnect_0:sram_controller_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_write;         // mm_interconnect_0:sram_controller_avalon_sram_slave_write -> sram_controller:write
	wire  [15:0] mm_interconnect_0_sram_controller_avalon_sram_slave_writedata;     // mm_interconnect_0:sram_controller_avalon_sram_slave_writedata -> sram_controller:writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata;      // pixel_buffer:slave_readdata -> mm_interconnect_0:pixel_buffer_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_address;       // mm_interconnect_0:pixel_buffer_avalon_control_slave_address -> pixel_buffer:slave_address
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_read;          // mm_interconnect_0:pixel_buffer_avalon_control_slave_read -> pixel_buffer:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable;    // mm_interconnect_0:pixel_buffer_avalon_control_slave_byteenable -> pixel_buffer:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_write;         // mm_interconnect_0:pixel_buffer_avalon_control_slave_write -> pixel_buffer:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata;     // mm_interconnect_0:pixel_buffer_avalon_control_slave_writedata -> pixel_buffer:slave_writedata
	wire  [31:0] mm_interconnect_0_resample_24bit_avalon_rgb_slave_readdata;        // resample_24bit:slave_readdata -> mm_interconnect_0:resample_24bit_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_resample_24bit_avalon_rgb_slave_read;            // mm_interconnect_0:resample_24bit_avalon_rgb_slave_read -> resample_24bit:slave_read
	wire  [31:0] mm_interconnect_0_vga_resample_avalon_rgb_slave_readdata;          // vga_resample:slave_readdata -> mm_interconnect_0:vga_resample_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_vga_resample_avalon_rgb_slave_read;              // mm_interconnect_0:vga_resample_avalon_rgb_slave_read -> vga_resample:slave_read
	wire  [31:0] mm_interconnect_0_resample_1bit_avalon_rgb_slave_readdata;         // resample_1bit:slave_readdata -> mm_interconnect_0:resample_1bit_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_resample_1bit_avalon_rgb_slave_read;             // mm_interconnect_0:resample_1bit_avalon_rgb_slave_read -> resample_1bit:slave_read
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;                   // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;                // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;                // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;                    // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;                       // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;                 // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;                      // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;                  // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                     // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_readdata;                       // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                        // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [1:0] mm_interconnect_0_onchip_memory_s1_byteenable;                     // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                          // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_writedata;                      // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                          // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         irq_mapper_receiver0_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_irq_irq;                                                      // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [dual_clock_buffer:reset_stream_in, edge_detector:reset, grayscale_converter:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:pixel_buffer_reset_reset_bridge_in_reset_reset, nios:reset_n, onchip_memory:reset, pixel_buffer:reset, pll_vga:ref_reset_reset, resample_1bit:reset, resample_24bit:reset, rst_translator:in_reset, scaler:reset, sram_controller:reset, vga_resample:reset]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [nios:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                                    // nios:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> dual_clock_buffer:reset_stream_out
	wire         pll_vga_reset_source_reset;                                        // pll_vga:reset_source_reset -> [rst_controller_001:reset_in2, rst_controller_002:reset_in0]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> vga_controller:reset

	IntegracaoPlatformDesigner_dual_clock_buffer dual_clock_buffer (
		.clk_stream_in            (clk_clk),                                                 //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                          //         reset_stream_in.reset
		.clk_stream_out           (pll_vga_vga_clk_clk),                                     //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                      //        reset_stream_out.reset
		.stream_in_ready          (scaler_avalon_scaler_source_ready),                       //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (scaler_avalon_scaler_source_startofpacket),               //                        .startofpacket
		.stream_in_endofpacket    (scaler_avalon_scaler_source_endofpacket),                 //                        .endofpacket
		.stream_in_valid          (scaler_avalon_scaler_source_valid),                       //                        .valid
		.stream_in_data           (scaler_avalon_scaler_source_data),                        //                        .data
		.stream_out_ready         (dual_clock_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	IntegracaoPlatformDesigner_edge_detector edge_detector (
		.clk               (clk_clk),                                                  //                          clk.clk
		.reset             (rst_controller_reset_out_reset),                           //                        reset.reset
		.in_data           (grayscale_converter_avalon_csc_source_data),               //   avalon_edge_detection_sink.data
		.in_startofpacket  (grayscale_converter_avalon_csc_source_startofpacket),      //                             .startofpacket
		.in_endofpacket    (grayscale_converter_avalon_csc_source_endofpacket),        //                             .endofpacket
		.in_valid          (grayscale_converter_avalon_csc_source_valid),              //                             .valid
		.in_ready          (grayscale_converter_avalon_csc_source_ready),              //                             .ready
		.out_ready         (edge_detector_avalon_edge_detection_source_ready),         // avalon_edge_detection_source.ready
		.out_data          (edge_detector_avalon_edge_detection_source_data),          //                             .data
		.out_startofpacket (edge_detector_avalon_edge_detection_source_startofpacket), //                             .startofpacket
		.out_endofpacket   (edge_detector_avalon_edge_detection_source_endofpacket),   //                             .endofpacket
		.out_valid         (edge_detector_avalon_edge_detection_source_valid)          //                             .valid
	);

	IntegracaoPlatformDesigner_grayscale_converter grayscale_converter (
		.clk                      (clk_clk),                                             //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //             reset.reset
		.stream_in_startofpacket  (resample_24bit_avalon_rgb_source_startofpacket),      //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (resample_24bit_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_in_valid          (resample_24bit_avalon_rgb_source_valid),              //                  .valid
		.stream_in_ready          (resample_24bit_avalon_rgb_source_ready),              //                  .ready
		.stream_in_data           (resample_24bit_avalon_rgb_source_data),               //                  .data
		.stream_out_ready         (grayscale_converter_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (grayscale_converter_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (grayscale_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (grayscale_converter_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (grayscale_converter_avalon_csc_source_data)           //                  .data
	);

	IntegracaoPlatformDesigner_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	IntegracaoPlatformDesigner_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	IntegracaoPlatformDesigner_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	IntegracaoPlatformDesigner_pixel_buffer pixel_buffer (
		.clk                  (clk_clk),                                                        //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (pixel_buffer_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_avalon_pixel_source_data)                           //                        .data
	);

	IntegracaoPlatformDesigner_pll_vga pll_vga (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (pll_vga_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset (pll_vga_reset_source_reset)      // reset_source.reset
	);

	IntegracaoPlatformDesigner_resample_1bit resample_1bit (
		.clk                      (clk_clk),                                                   //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                            //             reset.reset
		.stream_in_startofpacket  (edge_detector_avalon_edge_detection_source_startofpacket),  //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (edge_detector_avalon_edge_detection_source_endofpacket),    //                  .endofpacket
		.stream_in_valid          (edge_detector_avalon_edge_detection_source_valid),          //                  .valid
		.stream_in_ready          (edge_detector_avalon_edge_detection_source_ready),          //                  .ready
		.stream_in_data           (edge_detector_avalon_edge_detection_source_data),           //                  .data
		.slave_read               (mm_interconnect_0_resample_1bit_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_resample_1bit_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (resample_1bit_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (resample_1bit_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (resample_1bit_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (resample_1bit_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (resample_1bit_avalon_rgb_source_data)                       //                  .data
	);

	IntegracaoPlatformDesigner_resample_24bit resample_24bit (
		.clk                      (clk_clk),                                                    //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                             //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_avalon_pixel_source_startofpacket),             //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_avalon_pixel_source_endofpacket),               //                  .endofpacket
		.stream_in_valid          (pixel_buffer_avalon_pixel_source_valid),                     //                  .valid
		.stream_in_ready          (pixel_buffer_avalon_pixel_source_ready),                     //                  .ready
		.stream_in_data           (pixel_buffer_avalon_pixel_source_data),                      //                  .data
		.slave_read               (mm_interconnect_0_resample_24bit_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_resample_24bit_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (resample_24bit_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (resample_24bit_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (resample_24bit_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (resample_24bit_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (resample_24bit_avalon_rgb_source_data)                       //                  .data
	);

	IntegracaoPlatformDesigner_scaler scaler (
		.clk                      (clk_clk),                                      //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),               //                reset.reset
		.stream_in_startofpacket  (vga_resample_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (vga_resample_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (vga_resample_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (vga_resample_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (vga_resample_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),            // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),    //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),      //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),            //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data)              //                     .data
	);

	altera_external_memory_bfm #(
		.USE_CHIPSELECT           (1),
		.USE_WRITE                (1),
		.USE_READ                 (0),
		.USE_OUTPUTENABLE         (1),
		.USE_BEGINTRANSFER        (0),
		.ACTIVE_LOW_BYTEENABLE    (1),
		.ACTIVE_LOW_CHIPSELECT    (1),
		.ACTIVE_LOW_WRITE         (1),
		.ACTIVE_LOW_READ          (0),
		.ACTIVE_LOW_OUTPUTENABLE  (1),
		.ACTIVE_LOW_BEGINTRANSFER (0),
		.ACTIVE_LOW_RESET         (0),
		.CDT_ADDRESS_W            (20),
		.CDT_SYMBOL_W             (8),
		.CDT_NUMSYMBOLS           (2),
		.INIT_FILE                ("altera_external_memory_bfm.hex"),
		.CDT_READ_LATENCY         (2),
		.VHDL_ID                  (0)
	) sram (
		.clk               (clk_clk),                       //     clk.clk
		.cdt_write         (sram_conduit_cdt_write),        // conduit.cdt_write
		.cdt_chipselect    (sram_conduit_cdt_chipselect),   //        .cdt_chipselect
		.cdt_outputenable  (sram_conduit_cdt_outputenable), //        .cdt_outputenable
		.cdt_address       (sram_conduit_cdt_address),      //        .cdt_address
		.cdt_data_io       (sram_conduit_cdt_data_io),      //        .cdt_data_io
		.cdt_byteenable    (sram_conduit_cdt_byteenable),   //        .cdt_byteenable
		.cdt_read          (1'b0),                          // (terminated)
		.cdt_begintransfer (1'b0),                          // (terminated)
		.cdt_reset         (1'b0)                           // (terminated)
	);

	IntegracaoPlatformDesigner_sram_controller sram_controller (
		.clk           (clk_clk),                                                           //                clk.clk
		.reset         (rst_controller_reset_out_reset),                                    //              reset.reset
		.SRAM_DQ       (sram_controller_conduit_DQ),                                        // external_interface.export
		.SRAM_ADDR     (sram_controller_conduit_ADDR),                                      //                   .export
		.SRAM_LB_N     (sram_controller_conduit_LB_N),                                      //                   .export
		.SRAM_UB_N     (sram_controller_conduit_UB_N),                                      //                   .export
		.SRAM_CE_N     (sram_controller_conduit_CE_N),                                      //                   .export
		.SRAM_OE_N     (sram_controller_conduit_OE_N),                                      //                   .export
		.SRAM_WE_N     (sram_controller_conduit_WE_N),                                      //                   .export
		.address       (mm_interconnect_0_sram_controller_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_controller_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_controller_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_controller_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_controller_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	IntegracaoPlatformDesigner_vga_controller vga_controller (
		.clk           (pll_vga_vga_clk_clk),                                     //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                      //              reset.reset
		.data          (dual_clock_buffer_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_buffer_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_buffer_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_conduit_CLK),                                         // external_interface.export
		.VGA_HS        (vga_conduit_HS),                                          //                   .export
		.VGA_VS        (vga_conduit_VS),                                          //                   .export
		.VGA_BLANK     (vga_conduit_BLANK),                                       //                   .export
		.VGA_SYNC      (vga_conduit_SYNC),                                        //                   .export
		.VGA_R         (vga_conduit_R),                                           //                   .export
		.VGA_G         (vga_conduit_G),                                           //                   .export
		.VGA_B         (vga_conduit_B)                                            //                   .export
	);

	IntegracaoPlatformDesigner_vga_resample vga_resample (
		.clk                      (clk_clk),                                                  //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                           //             reset.reset
		.stream_in_startofpacket  (resample_1bit_avalon_rgb_source_startofpacket),            //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (resample_1bit_avalon_rgb_source_endofpacket),              //                  .endofpacket
		.stream_in_valid          (resample_1bit_avalon_rgb_source_valid),                    //                  .valid
		.stream_in_ready          (resample_1bit_avalon_rgb_source_ready),                    //                  .ready
		.stream_in_data           (resample_1bit_avalon_rgb_source_data),                     //                  .data
		.slave_read               (mm_interconnect_0_vga_resample_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_vga_resample_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (vga_resample_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (vga_resample_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (vga_resample_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (vga_resample_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (vga_resample_avalon_rgb_source_data)                       //                  .data
	);

	IntegracaoPlatformDesigner_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                                           //                                  clk_clk.clk
		.pixel_buffer_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                    // pixel_buffer_reset_reset_bridge_in_reset.reset
		.nios_data_master_address                           (nios_data_master_address),                                          //                         nios_data_master.address
		.nios_data_master_waitrequest                       (nios_data_master_waitrequest),                                      //                                         .waitrequest
		.nios_data_master_byteenable                        (nios_data_master_byteenable),                                       //                                         .byteenable
		.nios_data_master_read                              (nios_data_master_read),                                             //                                         .read
		.nios_data_master_readdata                          (nios_data_master_readdata),                                         //                                         .readdata
		.nios_data_master_write                             (nios_data_master_write),                                            //                                         .write
		.nios_data_master_writedata                         (nios_data_master_writedata),                                        //                                         .writedata
		.nios_data_master_debugaccess                       (nios_data_master_debugaccess),                                      //                                         .debugaccess
		.nios_instruction_master_address                    (nios_instruction_master_address),                                   //                  nios_instruction_master.address
		.nios_instruction_master_waitrequest                (nios_instruction_master_waitrequest),                               //                                         .waitrequest
		.nios_instruction_master_read                       (nios_instruction_master_read),                                      //                                         .read
		.nios_instruction_master_readdata                   (nios_instruction_master_readdata),                                  //                                         .readdata
		.pixel_buffer_avalon_pixel_dma_master_address       (pixel_buffer_avalon_pixel_dma_master_address),                      //     pixel_buffer_avalon_pixel_dma_master.address
		.pixel_buffer_avalon_pixel_dma_master_waitrequest   (pixel_buffer_avalon_pixel_dma_master_waitrequest),                  //                                         .waitrequest
		.pixel_buffer_avalon_pixel_dma_master_read          (pixel_buffer_avalon_pixel_dma_master_read),                         //                                         .read
		.pixel_buffer_avalon_pixel_dma_master_readdata      (pixel_buffer_avalon_pixel_dma_master_readdata),                     //                                         .readdata
		.pixel_buffer_avalon_pixel_dma_master_readdatavalid (pixel_buffer_avalon_pixel_dma_master_readdatavalid),                //                                         .readdatavalid
		.pixel_buffer_avalon_pixel_dma_master_lock          (pixel_buffer_avalon_pixel_dma_master_lock),                         //                                         .lock
		.jtag_uart_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),             //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),               //                                         .write
		.jtag_uart_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),            //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),           //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),         //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),          //                                         .chipselect
		.nios_debug_mem_slave_address                       (mm_interconnect_0_nios_debug_mem_slave_address),                    //                     nios_debug_mem_slave.address
		.nios_debug_mem_slave_write                         (mm_interconnect_0_nios_debug_mem_slave_write),                      //                                         .write
		.nios_debug_mem_slave_read                          (mm_interconnect_0_nios_debug_mem_slave_read),                       //                                         .read
		.nios_debug_mem_slave_readdata                      (mm_interconnect_0_nios_debug_mem_slave_readdata),                   //                                         .readdata
		.nios_debug_mem_slave_writedata                     (mm_interconnect_0_nios_debug_mem_slave_writedata),                  //                                         .writedata
		.nios_debug_mem_slave_byteenable                    (mm_interconnect_0_nios_debug_mem_slave_byteenable),                 //                                         .byteenable
		.nios_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios_debug_mem_slave_waitrequest),                //                                         .waitrequest
		.nios_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios_debug_mem_slave_debugaccess),                //                                         .debugaccess
		.onchip_memory_s1_address                           (mm_interconnect_0_onchip_memory_s1_address),                        //                         onchip_memory_s1.address
		.onchip_memory_s1_write                             (mm_interconnect_0_onchip_memory_s1_write),                          //                                         .write
		.onchip_memory_s1_readdata                          (mm_interconnect_0_onchip_memory_s1_readdata),                       //                                         .readdata
		.onchip_memory_s1_writedata                         (mm_interconnect_0_onchip_memory_s1_writedata),                      //                                         .writedata
		.onchip_memory_s1_byteenable                        (mm_interconnect_0_onchip_memory_s1_byteenable),                     //                                         .byteenable
		.onchip_memory_s1_chipselect                        (mm_interconnect_0_onchip_memory_s1_chipselect),                     //                                         .chipselect
		.onchip_memory_s1_clken                             (mm_interconnect_0_onchip_memory_s1_clken),                          //                                         .clken
		.pixel_buffer_avalon_control_slave_address          (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),       //        pixel_buffer_avalon_control_slave.address
		.pixel_buffer_avalon_control_slave_write            (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),         //                                         .write
		.pixel_buffer_avalon_control_slave_read             (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),          //                                         .read
		.pixel_buffer_avalon_control_slave_readdata         (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),      //                                         .readdata
		.pixel_buffer_avalon_control_slave_writedata        (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),     //                                         .writedata
		.pixel_buffer_avalon_control_slave_byteenable       (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable),    //                                         .byteenable
		.resample_1bit_avalon_rgb_slave_read                (mm_interconnect_0_resample_1bit_avalon_rgb_slave_read),             //           resample_1bit_avalon_rgb_slave.read
		.resample_1bit_avalon_rgb_slave_readdata            (mm_interconnect_0_resample_1bit_avalon_rgb_slave_readdata),         //                                         .readdata
		.resample_24bit_avalon_rgb_slave_read               (mm_interconnect_0_resample_24bit_avalon_rgb_slave_read),            //          resample_24bit_avalon_rgb_slave.read
		.resample_24bit_avalon_rgb_slave_readdata           (mm_interconnect_0_resample_24bit_avalon_rgb_slave_readdata),        //                                         .readdata
		.sram_controller_avalon_sram_slave_address          (mm_interconnect_0_sram_controller_avalon_sram_slave_address),       //        sram_controller_avalon_sram_slave.address
		.sram_controller_avalon_sram_slave_write            (mm_interconnect_0_sram_controller_avalon_sram_slave_write),         //                                         .write
		.sram_controller_avalon_sram_slave_read             (mm_interconnect_0_sram_controller_avalon_sram_slave_read),          //                                         .read
		.sram_controller_avalon_sram_slave_readdata         (mm_interconnect_0_sram_controller_avalon_sram_slave_readdata),      //                                         .readdata
		.sram_controller_avalon_sram_slave_writedata        (mm_interconnect_0_sram_controller_avalon_sram_slave_writedata),     //                                         .writedata
		.sram_controller_avalon_sram_slave_byteenable       (mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable),    //                                         .byteenable
		.sram_controller_avalon_sram_slave_readdatavalid    (mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid), //                                         .readdatavalid
		.vga_resample_avalon_rgb_slave_read                 (mm_interconnect_0_vga_resample_avalon_rgb_slave_read),              //            vga_resample_avalon_rgb_slave.read
		.vga_resample_avalon_rgb_slave_readdata             (mm_interconnect_0_vga_resample_avalon_rgb_slave_readdata)           //                                         .readdata
	);

	IntegracaoPlatformDesigner_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.reset_in2      (pll_vga_reset_source_reset),         // reset_in2.reset
		.clk            (pll_vga_vga_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (pll_vga_reset_source_reset),         // reset_in0.reset
		.clk            (pll_vga_vga_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
