// IntegracaoPlatformDesigner_tb.v

// Generated using ACDS version 20.1 720

`timescale 1 ns / 1 ns
module IntegracaoPlatformDesigner_tb (
	);

    integer      arquivo;
	wire         integracaoplatformdesigner_inst_clk_bfm_clk_clk;                           // IntegracaoPlatformDesigner_inst_clk_bfm:clk -> [IntegracaoPlatformDesigner_inst:clk_clk, IntegracaoPlatformDesigner_inst_reset_bfm:clk]
	wire  [19:0] integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_address;      // IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_address -> IntegracaoPlatformDesigner_inst:sram_conduit_cdt_address
	wire   [0:0] integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_outputenable; // IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_outputenable -> IntegracaoPlatformDesigner_inst:sram_conduit_cdt_outputenable
	wire  [15:0] integracaoplatformdesigner_inst_sram_conduit_cdt_data_io;                  // [] -> [IntegracaoPlatformDesigner_inst:sram_conduit_cdt_data_io, IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_data_io]
	wire   [0:0] integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_chipselect;   // IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_chipselect -> IntegracaoPlatformDesigner_inst:sram_conduit_cdt_chipselect
	wire   [0:0] integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_write;        // IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_write -> IntegracaoPlatformDesigner_inst:sram_conduit_cdt_write
	wire   [1:0] integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_byteenable;   // IntegracaoPlatformDesigner_inst_sram_conduit_bfm:sig_cdt_byteenable -> IntegracaoPlatformDesigner_inst:sram_conduit_cdt_byteenable
	wire         integracaoplatformdesigner_inst_sram_controller_conduit_oe_n;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_OE_N -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_OE_N
	wire         integracaoplatformdesigner_inst_sram_controller_conduit_we_n;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_WE_N -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_WE_N
	wire         integracaoplatformdesigner_inst_sram_controller_conduit_lb_n;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_LB_N -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_LB_N
	wire         integracaoplatformdesigner_inst_sram_controller_conduit_ub_n;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_UB_N -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_UB_N
	wire  [15:0] integracaoplatformdesigner_inst_sram_controller_conduit_dq;                // [] -> [IntegracaoPlatformDesigner_inst:sram_controller_conduit_DQ, IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_DQ]
	wire         integracaoplatformdesigner_inst_sram_controller_conduit_ce_n;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_CE_N -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_CE_N
	wire  [19:0] integracaoplatformdesigner_inst_sram_controller_conduit_addr;              // IntegracaoPlatformDesigner_inst:sram_controller_conduit_ADDR -> IntegracaoPlatformDesigner_inst_sram_controller_conduit_bfm:sig_ADDR
	wire         integracaoplatformdesigner_inst_vga_conduit_blank;                         // IntegracaoPlatformDesigner_inst:vga_conduit_BLANK -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_BLANK
	wire   [7:0] integracaoplatformdesigner_inst_vga_conduit_b;                             // IntegracaoPlatformDesigner_inst:vga_conduit_B -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_B
	wire   [7:0] integracaoplatformdesigner_inst_vga_conduit_r;                             // IntegracaoPlatformDesigner_inst:vga_conduit_R -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_R
	wire         integracaoplatformdesigner_inst_vga_conduit_clk;                           // IntegracaoPlatformDesigner_inst:vga_conduit_CLK -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_CLK
	wire   [7:0] integracaoplatformdesigner_inst_vga_conduit_g;                             // IntegracaoPlatformDesigner_inst:vga_conduit_G -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_G
	wire         integracaoplatformdesigner_inst_vga_conduit_hs;                            // IntegracaoPlatformDesigner_inst:vga_conduit_HS -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_HS
	wire         integracaoplatformdesigner_inst_vga_conduit_sync;                          // IntegracaoPlatformDesigner_inst:vga_conduit_SYNC -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_SYNC
	wire         integracaoplatformdesigner_inst_vga_conduit_vs;                            // IntegracaoPlatformDesigner_inst:vga_conduit_VS -> IntegracaoPlatformDesigner_inst_vga_conduit_bfm:sig_VS
	wire         integracaoplatformdesigner_inst_reset_bfm_reset_reset;                     // IntegracaoPlatformDesigner_inst_reset_bfm:reset -> IntegracaoPlatformDesigner_inst:reset_reset_n

	IntegracaoPlatformDesigner integracaoplatformdesigner_inst (
		.clk_clk                       (integracaoplatformdesigner_inst_clk_bfm_clk_clk),                           //                     clk.clk
		.reset_reset_n                 (integracaoplatformdesigner_inst_reset_bfm_reset_reset),                     //                   reset.reset_n
		.sram_conduit_cdt_write        (integracaoplatformdesigner_inst_sram_controller_conduit_we_n),        //            sram_conduit.cdt_write
		.sram_conduit_cdt_chipselect   (integracaoplatformdesigner_inst_sram_controller_conduit_ce_n),   //                        .cdt_chipselect
		.sram_conduit_cdt_outputenable (integracaoplatformdesigner_inst_sram_controller_conduit_oe_n), //                        .cdt_outputenable
		.sram_conduit_cdt_address      (integracaoplatformdesigner_inst_sram_controller_conduit_addr),      //                        .cdt_address
		.sram_conduit_cdt_data_io      (integracaoplatformdesigner_inst_sram_controller_conduit_dq),                  //                        .cdt_data_io
		.sram_conduit_cdt_byteenable   ({integracaoplatformdesigner_inst_sram_controller_conduit_ub_n, integracaoplatformdesigner_inst_sram_controller_conduit_lb_n}),   //                        .cdt_byteenable
		.sram_controller_conduit_DQ    (integracaoplatformdesigner_inst_sram_controller_conduit_dq),                // sram_controller_conduit.DQ
		.sram_controller_conduit_ADDR  (integracaoplatformdesigner_inst_sram_controller_conduit_addr),              //                        .ADDR
		.sram_controller_conduit_LB_N  (integracaoplatformdesigner_inst_sram_controller_conduit_lb_n),              //                        .LB_N
		.sram_controller_conduit_UB_N  (integracaoplatformdesigner_inst_sram_controller_conduit_ub_n),              //                        .UB_N
		.sram_controller_conduit_CE_N  (integracaoplatformdesigner_inst_sram_controller_conduit_ce_n),              //                        .CE_N
		.sram_controller_conduit_OE_N  (integracaoplatformdesigner_inst_sram_controller_conduit_oe_n),              //                        .OE_N
		.sram_controller_conduit_WE_N  (integracaoplatformdesigner_inst_sram_controller_conduit_we_n),              //                        .WE_N
		.vga_conduit_CLK               (integracaoplatformdesigner_inst_vga_conduit_clk),                           //             vga_conduit.CLK
		.vga_conduit_HS                (integracaoplatformdesigner_inst_vga_conduit_hs),                            //                        .HS
		.vga_conduit_VS                (integracaoplatformdesigner_inst_vga_conduit_vs),                            //                        .VS
		.vga_conduit_BLANK             (integracaoplatformdesigner_inst_vga_conduit_blank),                         //                        .BLANK
		.vga_conduit_SYNC              (integracaoplatformdesigner_inst_vga_conduit_sync),                          //                        .SYNC
		.vga_conduit_R                 (integracaoplatformdesigner_inst_vga_conduit_r),                             //                        .R
		.vga_conduit_G                 (integracaoplatformdesigner_inst_vga_conduit_g),                             //                        .G
		.vga_conduit_B                 (integracaoplatformdesigner_inst_vga_conduit_b)                              //                        .B
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) integracaoplatformdesigner_inst_clk_bfm (
		.clk (integracaoplatformdesigner_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) integracaoplatformdesigner_inst_reset_bfm (
		.reset (integracaoplatformdesigner_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (integracaoplatformdesigner_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm integracaoplatformdesigner_inst_sram_conduit_bfm (
		.sig_cdt_address      (integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_address),      // conduit.cdt_address
		.sig_cdt_byteenable   (integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_byteenable),   //        .cdt_byteenable
		.sig_cdt_chipselect   (integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_chipselect),   //        .cdt_chipselect
		.sig_cdt_data_io      (integracaoplatformdesigner_inst_sram_conduit_cdt_data_io),                  //        .cdt_data_io
		.sig_cdt_outputenable (integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_outputenable), //        .cdt_outputenable
		.sig_cdt_write        (integracaoplatformdesigner_inst_sram_conduit_bfm_conduit_cdt_write)         //        .cdt_write
	);

	altera_conduit_bfm_0002 integracaoplatformdesigner_inst_sram_controller_conduit_bfm (
		.sig_ADDR (integracaoplatformdesigner_inst_sram_controller_conduit_addr), // conduit.ADDR
		.sig_CE_N (integracaoplatformdesigner_inst_sram_controller_conduit_ce_n), //        .CE_N
		.sig_DQ   (integracaoplatformdesigner_inst_sram_controller_conduit_dq),   //        .DQ
		.sig_LB_N (integracaoplatformdesigner_inst_sram_controller_conduit_lb_n), //        .LB_N
		.sig_OE_N (integracaoplatformdesigner_inst_sram_controller_conduit_oe_n), //        .OE_N
		.sig_UB_N (integracaoplatformdesigner_inst_sram_controller_conduit_ub_n), //        .UB_N
		.sig_WE_N (integracaoplatformdesigner_inst_sram_controller_conduit_we_n)  //        .WE_N
	);

	altera_conduit_bfm_0003 integracaoplatformdesigner_inst_vga_conduit_bfm (
		.sig_B     (integracaoplatformdesigner_inst_vga_conduit_b),     // conduit.B
		.sig_BLANK (integracaoplatformdesigner_inst_vga_conduit_blank), //        .BLANK
		.sig_CLK   (integracaoplatformdesigner_inst_vga_conduit_clk),   //        .CLK
		.sig_G     (integracaoplatformdesigner_inst_vga_conduit_g),     //        .G
		.sig_HS    (integracaoplatformdesigner_inst_vga_conduit_hs),    //        .HS
		.sig_R     (integracaoplatformdesigner_inst_vga_conduit_r),     //        .R
		.sig_SYNC  (integracaoplatformdesigner_inst_vga_conduit_sync),  //        .SYNC
		.sig_VS    (integracaoplatformdesigner_inst_vga_conduit_vs)     //        .VS
	);

	initial begin
        arquivo = $fopen("imageoutputnios.txt", "w");         
	end

	always @ (posedge integracaoplatformdesigner_inst_vga_conduit_clk) begin
		if ($time > 16700000 && integracaoplatformdesigner_inst_vga_conduit_vs == 0) begin // segundo frame
		//if ($time > 340 && integracaoplatformdesigner_inst_vga_conduit_vs == 0) begin // primeiro frame
			$fclose(arquivo);
		end
		else begin
			if($time > 16700000 && integracaoplatformdesigner_inst_vga_conduit_blank != 0) begin // segundo frame
			//if($time > 340 && integracaoplatformdesigner_inst_vga_conduit_blank != 0) begin // primeiro frame
				$fwrite(arquivo,"00000000%b%b%b\n", integracaoplatformdesigner_inst_vga_conduit_r, integracaoplatformdesigner_inst_vga_conduit_g, integracaoplatformdesigner_inst_vga_conduit_b);
			end
		end
	end

endmodule
